//////////////////////////////////////////////////////////////////////////////////
// Company:         University of Duisburg-Essen, Intelligent Embedded Systems Lab
// Engineer:        AE
// 
// Create Date:     13.01.2025 23:07:45
// Copied on: 	    {$date_copy_created}
// Module Name:     SKELETON_DNN
// Target Devices:  FPGA
// Tool Versions:   1v0
// Description:     Skeleton for testing Deep Learning models, generated by elasticAI.creator on device
// Dependencies:    None
//
// State: 	        Works! (System Test done: 16.01.2025)
// Improvements:    None
// Parameters:      BITWIDTH_IN 	--> Bitwidth of input data
//                  BITWIDTH_SYS 	--> Bitwidth of data bus on device
//                  BITWIDTH_HEAD	--> Bitwidth of metadata (skeleton properties)
//					ADR_WIDTH 		--> Bitwidth of adress range
//////////////////////////////////////////////////////////////////////////////////


module SKELETON_NN#(
	parameter BITWIDTH_IN = 5'd8,
    parameter BITWIDTH_SYS = 5'd16,
    parameter BITWIDTH_HEAD = 6'd32,
	parameter ADR_WIDTH = 6'd6
)(
    input wire CLK,
    input wire nRST,
    input wire EN,
    input wire RnW,
    input wire [ADR_WIDTH-'d1:0] ADR,
    input wire [BITWIDTH_SYS-'d1:0] DATA_IN,
    output wire [BITWIDTH_SYS-'d1:0] DATA_OUT,
    output wire [BITWIDTH_HEAD-'d7:0] DATA_HEAD,
	output wire DATA_VALID
);

localparam BITWIDTH_OFFSET = BITWIDTH_SYS - BITWIDTH_IN;
assign DATA_HEAD = {4'd7, 6'd5, 6'd3, BITWIDTH_IN[4:0], BITWIDTH_IN[4:0]};
assign DATA_OUT[0+:BITWIDTH_OFFSET] = 8'd0;

//If using skeleton from elasticAI.creator please include shift, otherwise software API does not work!
//Also include SEL in reset input
skeleton LinearDesign(
    .clock(CLK),
    .clk_hadamard(CLK),
    .reset(~(nRST && EN)),
    .busy(DATA_VALID),
    .wake_up(),
    .rd(RnW),
    .wr(~RnW),
    .data_in(DATA_IN[BITWIDTH_OFFSET+:BITWIDTH_IN]),
    .address_in({{('d16-ADR_WIDTH){1'd0}}, ADR}),    
    .data_out(DATA_OUT[BITWIDTH_OFFSET+:BITWIDTH_IN]),
    .debug()
);


endmodule
