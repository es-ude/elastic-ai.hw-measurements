module TEST_ENVIRONMENT#(
    parameter BITWIDTH_DATA = 16,
    parameter BITWIDTH_ADR = 6,
    parameter NUM_DUT = 4,
    parameter NUM_BITS_HEADER = 32,
    parameter UINT_DATATYPE = 1
)(
    input wire CLK,
    input wire RSTN,
    input wire START_FLAG,
    input wire [$clog2(NUM_DUT):0] SEL,
    input wire [BITWIDTH_ADR-'d1:0] ADR,
    input wire RnW,
    input wire [BITWIDTH_DATA-'d1:0] DATA_IN,
    output wire [BITWIDTH_DATA-'d1:0] DATA_OUT,
    output wire [NUM_BITS_HEADER-'d1:0] HEAD_INFO, 
    output wire RDY_FLAG
);

    localparam BITWIDTH_HEAD = NUM_BITS_HEADER - 'd6;
    //################## CONTROL LINES ################## 
    wire [BITWIDTH_DATA-'d1:0] dout [NUM_DUT:0];
    assign DATA_OUT = dout[SEL]; 

    wire [NUM_DUT:0] rdy_filt;
    assign RDY_FLAG = rdy_filt[SEL];
    
    //* This variable contains information about the module for read-in in Python 
    //  - NUM_DUTS (6-bits):        Total number of DUTs available in this function (automated added here)
    //  - DUT_TPYE (4-bits):        0 = Echo, 1 = Multiplier, 2 = Division, 3 = ROM, 4 = RAM, 5 = Filter, 6 = Processor, 7 = Skeleton (elasticAI.creator)
    //  - NUM_INPUTS (6-bits):      Number of used inputs
    //  - NUM_OUTPUTS (6-bits):     Number of used outputs
    //  - BITWIDTH_IN (5-bits):     Bitwidth of input data
    //  - BITWIDTH_OUT (5-bits):    Bitwidth of output data
    wire [NUM_BITS_HEADER-'d7:0] head_array [NUM_DUT:0];
    assign HEAD_INFO = {NUM_DUT[5:0], head_array[SEL]};

    // SEL == 'd0 will be skipped!
    assign dout[0] = 'd0123;
    assign head_array[0] = {4'd0, 6'd0, 6'd1, 5'd0, BITWIDTH_DATA[4:0]};
    assign rdy_filt[0] = 1'd0; 

    //################## List with DUT ################## 
    SKELETON_ECHO#(BITWIDTH_DATA, BITWIDTH_HEAD) DUT_01 (
        .CLK_SYS(CLK),
        .RSTN(RSTN),
        .EN(SEL == 'd1),
        .TRGG_START_CALC(START_FLAG),
        .DATA_IN(DATA_IN),
        .DATA_OUT(dout[1]),
        .DATA_HEAD(head_array[1]),
        .DATA_VALID(rdy_filt[1])
    );    
        
    SKELETON_ROM#('d16, BITWIDTH_DATA, BITWIDTH_HEAD) DUT_02 (
        .CLK_SYS(CLK),
        .RSTN(RSTN),
		.EN(SEL == 'd2),
		.TRGG_START_CALC(START_FLAG),
		.DATA_IN(DATA_IN),
		.DATA_OUT(dout[2]),
		.DATA_HEAD(head_array[2]),
		.RDY(rdy_filt[2])
    );  
    
    SKELETON_RAM#('d16, BITWIDTH_DATA, BITWIDTH_HEAD, BITWIDTH_ADR) DUT_03 (
        .CLK_SYS(CLK),
        .RSTN(RSTN),
		.EN(SEL == 'd3),
		.TRGG_START_CALC(START_FLAG),
		.RnW(RnW),
		.ADR(ADR),
		.DATA_IN(DATA_IN),
		.DATA_OUT(dout[3]),
		.DATA_HEAD(head_array[3]),
		.RDY(rdy_filt[3])    
    );

    SKELETON_MATH#(
        .BITWIDTH_IN('d8),
        .BITWIDTH_SYS(BITWIDTH_DATA),
        .BITWIDTH_HEAD(BITWIDTH_HEAD),
        .BITWIDTH_ADR(BITWIDTH_ADR)
    ) DUT_04 (
        .CLK_SYS(CLK),
        .RSTN(RSTN),
		.EN(SEL == 'd4),
		.TRGG_START_CALC(START_FLAG),
		.RnW(RnW),
		.ADR(ADR),
		.DATA_IN(DATA_IN),
		.DATA_OUT(dout[4]),
		.DATA_HEAD(head_array[4]),
		.RDY(rdy_filt[4])
    );
        
endmodule
